/***********************************************************************************************************************
 * Copyright (c) 2024 Virgil Dobjanschi dobjanschivirgil@gmail.com
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy of this software and associated
 * documentation files (the "Software"), to deal in the Software without restriction, including without limitation the
 * rights to use, copy, modify, merge, publish, distribute, sublicense, and/or sell copies of the Software, and to
 * permit persons to whom the Software is furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in all copies or substantial portions of
 * the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE
 * WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS
 * OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR
 * OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
 **********************************************************************************************************************/

/***********************************************************************************************************************
 * RAM driver module for an SDRAM featuring a wishbone interface.
 *
 * ULX3S uses the IS42S16160G-7 SDRAM a 16 Meg x 16 SDRAM (4 Meg x 16 x 4 banks)
 * Rows     :8192   A[12:0]
 * Columns  :512    A[8:0]
 * Banks    :4      BA[1:0]
 *
 * clk_i        -- The clock signal.
 * rst_i        -- Reset active high.
 * stb_i        -- The data transaction starts on the posedge of this signal.
 * cyc_i        -- This signal is asserted for the duration of a cycle.
 * sel_i        -- The number of bytes to read (1 -> 4'b0001, 2 -> 4'b0011, 3 -> 4'b0111 or 4 bytes -> 4'b1111).
 * we_i         -- 1 to write data, 0 to read.
 * addr_i       -- The address from where data is read/written.
 * data_i       -- The input data to write.
 * ack_o        -- The data request is complete on the posedge of this signal.
 * data_o       -- The data that was read.
 * device_clk_i -- The device clk generated by the PLL.
 * SDRAM wires  -- SDRAM signals.
 **********************************************************************************************************************/
`timescale 1ns / 1ns
`default_nettype none

module sdram #(parameter [31:0] CLK_PERIOD_NS = 20) (
    // Wishbone interface
    input logic clk_i,
    input logic rst_i,
    input logic stb_i,
    input logic cyc_i,
    input logic [3:0] sel_i,
    input logic we_i,
    input logic [23:0] addr_i,
    input logic [31:0] data_i,
    output logic ack_o,
    output logic [31:0] data_o,
    // The device clock is driving sdram_clk
    input logic device_clk_i,
    // SDRAM signals
    output logic sdram_clk,
    output logic sdram_cke,
    output logic sdram_csn,
    output logic sdram_wen,
    output logic sdram_rasn,
    output logic sdram_casn,
    output logic [12:0] sdram_a,
    output logic [1:0] sdram_ba,
    output logic [1:0] sdram_dqm,
    inout logic [15:0] sdram_d);

    /*
     * Name (Function)                                          CS# RAS#    CAS#    WE#     DQM     ADDR        DQ
     * COMMAND INHIBIT (NOP)                                    H   X       X       X       X       X           X
     * NO OPERATION (NOP)                                       L   H       H       H       X       X           X
     * ACTIVE (select bank and activate row)                    L   L       H       H       X       Bank/row    X
     * READ (select bank and column, and start READ burst)      L   H       L       H       L/H     Bank/col    X
     * WRITE (select bank and column, and start WRITE burst)    L   H       L       L       L/H     Bank/col    Valid
     * BURST TERMINATE                                          L   H       H       L       X       X           Active
     * PRECHARGE (Deactivate row in bank or banks)              L   L       H       L       X       Code        X
     * AUTO REFRESH or SELF REFRESH                             L   L       L       H       X       X           X
     * LOAD MODE REGISTER                                       L   L       L       L       X       Op-code     X
     * Write enable/output enable                               X   X       X       X       L       X           Active
     * Write inhibit/output High-Z                              X   X       X       X       H       X           High-Z
     */

    /*
     * The NO OPERATION (NOP) command is used to perform a NOP to the selected device (CS# is LOW).
     * This prevents unwanted commands from being registered during idle or wait states.
     * Operations already in progress are not affected.
     */
    localparam [3:0] SDRAM_CMD_NOP = 4'b0111;
    /*
     * The ACTIVE command is used to activate a row in a particular bank for a subsequent access.
     * The value on the BA0, BA1 inputs selects the bank, and the address provided selects the row.
     * This row remains active for accesses until a PRECHARGE command is issued to that bank.
     * A PRECHARGE command must be issued before opening a different row in the same bank.
     */
    localparam [3:0] SDRAM_CMD_ACTIVE = 4'b0011;
    /*
     * The READ command is used to initiate a burst read access to an active row.
     * The values on the BA0 and BA1 inputs select the bank; the address provided selects the
     * starting column location.
     */
    localparam [3:0] SDRAM_CMD_READ = 4'b0101;
    /*
     * The WRITE command is used to initiate a burst write access to an active row.
     * The values on the BA0 and BA1 inputs select the bank; the address provided selects the
     * starting column location.
     */
    localparam [3:0] SDRAM_CMD_WRITE = 4'b0100;
    /*
     * The PRECHARGE command is used to deactivate the open row in a particular bank
     * or the open row in all banks.
     */
    localparam [3:0] SDRAM_CMD_PRECHARGE = 4'b0010;
    /*
     * AUTO REFRESH (CKE = H) is used during normal operation of the SDRAM and is analogous to
     * CAS#-BEFORE-RAS# (CBR) refresh in conventional DRAMs.
     * This command is nonpersistent, so it must be issued each time a refresh is required.
     */
    localparam [3:0] SDRAM_CMD_REFRESH = 4'b0001;
    /*
     * The mode registers are loaded via inputs A[n:0] (where An is the most significant address term), BA0, and BA1.
     */
    localparam [3:0] SDRAM_CMD_LOAD_MODE_REGISTER = 4'b0000;

    // The command to issue
    logic [3:0] sdram_cmd;
    assign {sdram_csn, sdram_rasn, sdram_casn, sdram_wen} = sdram_cmd;

    // Input/output 16-bit data bus
    logic [15:0] sdram_d_i, sdram_d_o;
    // .T = 0 -> sdram_d is output; .T = 1 -> sdram_d is input.
    TRELLIS_IO #(.DIR("BIDIR")) sdram_d_io[15:0] (.B(sdram_d), .I(sdram_d_o), .T(sdram_cmd != SDRAM_CMD_WRITE),
                            .O(sdram_d_i));

    // Drive the SDRAM clock with the clock generated by the PLL.
    assign sdram_clk = sdram_cke ? device_clk_i : 1'b0;

    // The wishbone ack_o is cleared as soon as stb_i is cleared.
    logic sync_ack_o = 1'b0;
    assign ack_o = sync_ack_o & stb_i;

    /* During reset bring CKE up sometime during this time interval (minimum 100μs) */
    localparam CKE_CLKS = 120000 / CLK_PERIOD_NS;
    /*
     * PRECHARGE command period: the bank(s) will be available for a subsequent row access a specified time (tRP)
     * after the PRECHARGE command is issued. tRP = minimum 15nS.
     */
    localparam TRP_CLKS = (20 / CLK_PERIOD_NS) + 1;
    /*
     * AUTO REFRESH commands can be issued in a burst at the minimum cycle rate (tRFC),
     * tRFC = minimum 60nS.
     */
    localparam TRFC_CLKS = (70 / CLK_PERIOD_NS) + 1;
    /*
     * The LOAD MODE REGISTER command can only be issued when all banks are idle and a subsequent executable
     * command cannot be issued until tMRD is met. tMRD = 14nS.
     */
    localparam TMRD_CLKS = 2;
    /*
     * After a row is opened with the ACTIVE command, a READ or WRITE command can be issued to that row,
     * subject to the tRCD specification. tRCD = minimum 20nS.
     */
    localparam TRCD_CLKS = (30 / CLK_PERIOD_NS) + 1;
    /*
     * Providing a distributed AUTO REFRESH command every 7.813μs (commercial and industrial) or
     * 1.953μs (automotive) will meet the refresh requirement and ensure that each row is refreshed.
     * This implementation uses 5μs.
     */
    localparam REFRESH_CLKS = 5000 / CLK_PERIOD_NS;

    // Reset machine states
    localparam STATE_RESET_BEGIN = 3'b000;
    localparam STATE_RESET_WAIT_HALF_CKE = 3'b001;
    localparam STATE_RESET_WAIT_CKE = 3'b010;
    localparam STATE_RESET_WAIT_TRP = 3'b011;
    localparam STATE_RESET_WAIT_TRFC = 3'b100;
    localparam STATE_RESET_WAIT_MRD = 3'b101;
    localparam STATE_RESET_END = 3'b110;
    // Reset state machine (rst_i == 1)
    logic [2:0] reset_state_m;

    // State machine for operation
    localparam STATE_RESET = 3'b000;
    localparam STATE_IDLE = 3'b001;
    localparam STATE_WAIT_TRCD = 3'b010;
    localparam STATE_ACTIVATED = 3'b011;
    localparam STATE_READ_PENDING = 3'b100;
    localparam STATE_PRECHARGE = 3'b101;
    localparam STATE_WAIT_TRP = 3'b110;
    localparam STATE_AUTO_REFRESH = 3'b111;
    // SDRAM controller state machine (rst_i == 0)
    logic [2:0] state_m;

    // Auto Refresh sub state machines
    localparam STATE_AR_START = 2'b00;
    localparam STATE_AR_WAIT_TRP = 2'b01;
    localparam STATE_AR_WAIT_TRFC = 2'b11;
    // Auto Refresh state machine (state_m == STATE_AUTO_REFRESH)
    logic [1:0] auto_refresh_state_m;

    // The default CAS latency is 2. cas_delay is used to shift a bit during read to implement the CAS latency.
    // Note: this code needs to wait an extra clock cycle to account for the delayed SDRAM clock.
    localparam CAS_DELAY = 2;
    logic [CAS_DELAY:0] cas_latency;

    logic [14:0] activated_row_bank;
    // This register is used to shift a bit during reset to indicate how many refresh cycles are performed.
    logic [1:0] reset_auto_refresh_count;
    // The following two bits are used to determine when a new transaction starts.
    logic prev_stb_cyc, transaction_start_q;
    logic reset_refresh_timer;
    logic next_word;
    logic [23:0] next_addr, active_addr;
    assign active_addr = next_word ? next_addr : addr_i;
    always_comb begin
        next_addr = addr_i + 1;
    end

    //==================================================================================================================
    // Precharge all banks task
    //==================================================================================================================
    task precharge_all_task;
        sdram_cmd <= SDRAM_CMD_PRECHARGE;
        sdram_ba  <= 0;
        // A10 = 1: all banks
        sdram_a   <= 13'b0_0100_0000_0000;
        sdram_dqm <= 2'b11;
    endtask

    //==================================================================================================================
    // The reset state machine
    //==================================================================================================================
    task reset_task;
        (* parallel_case, full_case *)
        case (reset_state_m)
            STATE_RESET_BEGIN: begin
                /*
                 * 1. Simultaneously apply power to V DD and V DDQ.
                 */
                sdram_dqm <= 2'b11;
                /*
                 * 2. Assert and hold CKE at a LVTTL logic LOW since all inputs and outputs are LVTTL-compatible.
                 */
                sdram_cke <= 1'b0;
                sdram_cmd <= SDRAM_CMD_NOP;
                /*
                 * 3. Provide stable CLOCK signal. Stable clock is defined as a signal cycling within
                 * timing constraints specified for the clock pin.
                 * Note that sdram_clk is enabled when sdram_cke is 1. See assign of sdram_clk above.
                 */
                set_timer_task(CKE_CLKS / 2);

                reset_state_m <= STATE_RESET_WAIT_HALF_CKE;
            end

            STATE_RESET_WAIT_HALF_CKE: begin
                if (timer_expired) begin
                    /*
                     * 5. Starting at some point during this 100μs period, bring CKE HIGH. Continuing at
                     * least through the end of this period, 1 or more COMMAND INHIBIT or NOP commands
                     * must be applied.
                     */
                    sdram_cke <= 1'b1;

                    set_timer_task(CKE_CLKS / 2);

                    reset_state_m <= STATE_RESET_WAIT_CKE;
                end
            end

            STATE_RESET_WAIT_CKE: begin
                /* 4. Wait at least 100μs prior to issuing any command other than a COMMAND INHIBIT/NOP.*/
                if (timer_expired) begin
                    /* 6. Perform a PRECHARGE ALL command.*/
                    precharge_all_task;

                    set_timer_task(TRP_CLKS);

                    reset_state_m <= STATE_RESET_WAIT_TRP;
                end
            end

            STATE_RESET_WAIT_TRP: begin
                /*
                 * 7. Wait at least tRP time; during this time NOPs or DESELECT commands must be given.
                 * All banks will complete their precharge, thereby placing the device in the all banks idle state.
                 */
                if (timer_expired) begin
                    /* 8. Issue an AUTO REFRESH command. */
                    sdram_cmd <= SDRAM_CMD_REFRESH;
                    /*
                     * Two cycles are required. We do 3, the one just started and then two more.
                     */
                    reset_auto_refresh_count <= 2'b10;

                    set_timer_task(TRFC_CLKS);

                    reset_state_m <= STATE_RESET_WAIT_TRFC;
                end else begin
                    sdram_cmd <= SDRAM_CMD_NOP;
                end
            end

            STATE_RESET_WAIT_TRFC: begin
                /*
                 * 9 & 11. Wait at least tRFC time, during which only NOPs or COMMAND INHIBIT commands are allowed.
                 */
                if (timer_expired) begin
                    if (reset_auto_refresh_count == 0) begin
                        /*
                         * 12. The SDRAM is now ready for mode register programming.
                         * Because the mode register will power up in an unknown state,
                         * it should be loaded with desired bit values prior to applying any operational
                         * command.
                         */
                        /*
                         * Using the LMR command, program the mode register.
                         * The mode register is programmed via the MODE REGISTER SET command with BA1 = 0,
                         * BA0 = 0 and retains the stored information until it is programmed again or the
                         * device loses power. Outputs should be High-Z  already before the LMR command is
                         * issued.
                         */
                        sdram_ba <= 2'b00;
                        /*
                         * Mode register bits M[2:0] specify the BL; We use BL = 1.
                         */
                        sdram_a[2:0] <= 3'b000;
                        /*
                         * M3 specifies the type of burst; Sequential is un use.
                         */
                        sdram_a[3] <= 1'b0;
                        /*
                         * M[6:4] specify the CL; We use 2 or 3.
                         */
                        sdram_a[6:4] <= CAS_DELAY;
                        /*
                         * M7 and M8 specify the operating mode. Standard Operation is enabled.
                         */
                        sdram_a[8:7] <= 2'b00;
                        /*
                         * M9 specifies the write burst mode; Single Location Access (disable burst) is enabled.
                         */
                        sdram_a[9] <= 1'b1;
                        /*
                         * and M10–Mn should be set to zero to ensure compatibility with future revisions.
                         * Mn + 1 and Mn + 2 should be set to zero to select the mode register.
                         */
                        sdram_a[12:10] <= 3'b000;

                        sdram_cmd <= SDRAM_CMD_LOAD_MODE_REGISTER;

                        set_timer_task(TMRD_CLKS);

                        reset_state_m <= STATE_RESET_WAIT_MRD;
                    end else begin
                        /* 10. Issue the next AUTO REFRESH command. */
                        sdram_cmd <= SDRAM_CMD_REFRESH;

                        reset_auto_refresh_count <= reset_auto_refresh_count - 1;

                        set_timer_task(TRFC_CLKS);
                        // Stay in this state machine
                    end
                end else begin
                    sdram_cmd <= SDRAM_CMD_NOP;
                end
            end

            STATE_RESET_WAIT_MRD: begin
                sdram_cmd <= SDRAM_CMD_NOP;

                if (timer_expired) begin
                    reset_state_m <= STATE_RESET_END;
                end
            end

            STATE_RESET_END: begin
`ifdef D_SDRAM
                $display($time, " SDRAM: SDRAM reset complete.");
`endif
                /* At this point the DRAM is ready for any valid command.*/
                activated_row_bank <= 0;
                state_m <= STATE_IDLE;
                next_word <= 1'b0;
            end

            default: begin
                // Invalid state machine
            end
        endcase
    endtask

    //==================================================================================================================
    // The multi-purpose timer task used by the main always block to start the timer.
    // Setting value to 0 will clear/cancel the timer. The main block needs to clear set_timer bit a clock after
    // executing the set_timer_task.
    //==================================================================================================================
    logic set_timer = 1'b0;
    logic [15:0] timer_set_value;  // The longest timer interval is for CKE_CLKS (12,000 cycles)

    task set_timer_task(input [15:0] value);
        timer_set_value <= value;
        set_timer <= 1'b1;
    endtask

    //==================================================================================================================
    // The multi-purpose timer implementation. Note that the timer is also used during reset.
    //==================================================================================================================
    logic timer_is_set = 1'b0;
    logic timer_expired = 1'b0;
    logic [15:0] timer_count;

    always @(posedge clk_i) begin

        timer_expired <= 1'b0;
        if (set_timer) begin
            (* parallel_case, full_case *)
            case (timer_set_value)
                0: begin
                    // Clear/cancel the timer
                    timer_is_set <= 1'b0;
                end

                1, 2: begin
                    // One clock cycle already passed and therefore the timer expired.
                    timer_is_set  <= 1'b0;
                    timer_expired <= 1'b1;
                end

                default: begin
                    timer_is_set <= 1'b1;
                    // One clock cycle already passed and one for one cycle late delivery of timer_expired.
                    timer_count  <= timer_set_value - 2;
                end
            endcase
        end else if (timer_is_set) begin
            if (timer_count == 1) begin
                timer_is_set  <= 1'b0;
                timer_expired <= 1'b1;
            end else begin
                timer_count <= timer_count - 1;
            end
        end
    end

    //==================================================================================================================
    // The refresh timer
    //==================================================================================================================
    logic refresh_expired;
    logic [10:0] refresh_counter;  // Maxiumum 2047 cycles (20μs @10ns CLK_PERIOD_NS)

    always @(posedge clk_i) begin
        if (rst_i) begin
            refresh_counter <= REFRESH_CLKS;
            refresh_expired <= 1'b0;
        end else begin
            if (reset_refresh_timer) begin
                refresh_counter <= REFRESH_CLKS;
                refresh_expired <= 1'b0;
            end else if (~|refresh_counter) begin
                refresh_expired <= 1'b1;
            end else begin
                refresh_counter <= refresh_counter - 1;
            end
        end
    end

    //==================================================================================================================
    // SDRAM controller
    //==================================================================================================================
    always @(posedge clk_i) begin
        if (rst_i) begin
            sync_ack_o <= 1'b0;
            transaction_start_q <= 1'b0;
            prev_stb_cyc <= 1'b0;

            cas_latency <= 0;

            reset_refresh_timer <= 1'b1;

            reset_state_m <= STATE_RESET_BEGIN;
            state_m <= STATE_RESET;
        end else begin
            // At the end of a transaction reset ack_o
            if (sync_ack_o) sync_ack_o <= stb_i;

            // Latch the request. We may not be able to service it right away.
            if (stb_i & cyc_i & ~ack_o & ~prev_stb_cyc) transaction_start_q <= 1'b1;
            prev_stb_cyc <= stb_i & cyc_i;

            reset_refresh_timer <= 1'b0;
            set_timer <= 1'b0;

            (* parallel_case, full_case *)
            case (state_m)
                STATE_RESET: begin
                    reset_task;
                end

                STATE_IDLE: begin
                    /*
                     * The address bits registered coincident with the ACTIVE command are used to select
                     * the bank and row to be accessed (BA[1:0] select the bank; A[12:0] select the row).
                     * The row remains active for accesses until a PRECHARGE command is issued to that bank.
                     * A PRECHARGE command must be issued before opening a different row in the same bank.
                     */
                    sdram_ba <= activated_row_bank[14:13];
                    sdram_a <= activated_row_bank[12:0];

                    // Activate the bank and the row
                    sdram_cmd <= SDRAM_CMD_ACTIVE;

                    /*
                     * After a row is opened with the ACTIVE command, a READ or WRITE command can be
                     * issued to that row, subject to the tRCD specification.
                     */
                    set_timer_task(TRCD_CLKS);

                    state_m <= STATE_WAIT_TRCD;
                end

                STATE_WAIT_TRCD: begin
                    sdram_cmd <= SDRAM_CMD_NOP;
                    if (timer_expired) begin
                        state_m <= STATE_ACTIVATED;
                    end
                end

                STATE_ACTIVATED: begin
                    if ((stb_i & cyc_i & ~ack_o & ~prev_stb_cyc) | transaction_start_q) begin
                        if (activated_row_bank == active_addr[23:9]) begin
                            // We started servicing this request
                            transaction_start_q <= 1'b0;
                            /*
                             * The READ/WRITE commands are used to initiate a burst read access to the active row.
                             * This is a read/write with the same bank and row as the last one. Just set the column.
                             * Auto precharge (A10) is disabled and therefore the row remains open for subsequent
                             * accesses.
                             */
                            sdram_a <= {4'b0000, active_addr[8:0]};
                            // DQM: Specify 0 for dqm[1] to get bites [15:8] and specify 0 for dqm[0] to get bits [7:0].
                            sdram_dqm <= ~sel_i[1:0];

                            if (we_i) begin
                                sdram_cmd <= SDRAM_CMD_WRITE;
                                if (sel_i[3]) begin
                                    if (next_word) begin
                                        sdram_d_o <= data_i[31:16];
                                        // The transaction is complete
                                        sync_ack_o <= 1'b1;
                                    end else begin
                                        sdram_d_o <= data_i[15:0];
                                        transaction_start_q <= 1'b1;
                                    end
                                    next_word <= ~next_word;
                                end else begin
                                    sdram_d_o <= data_i[15:0];
                                    // The transaction is complete
                                    sync_ack_o <= 1'b1;
                                end
                            end else begin
`ifdef D_SDRAM
                                $display($time,
                                    " SDRAM: STATE_ACTIVATED: Read: sel %h, @[%h]-> STATE_READ_PENDING (next word %h)",
                                            sel_i, active_addr, next_word);
`endif
                                // Read requests will complete when the bit is shifted left to the MSB of cas_latency.
                                cas_latency <= 1'b1;
                                sdram_cmd <= SDRAM_CMD_READ;
                                state_m <= STATE_READ_PENDING;
                            end
                        end else begin
                            activated_row_bank <= active_addr[23:9];
                            // Clear the bank and the row and activate the new bank and the new row.
                            sdram_cmd <= SDRAM_CMD_NOP;
                            state_m <= STATE_PRECHARGE;
`ifdef D_SDRAM
                            $display($time, " SDRAM: STATE_ACTIVATED: BR: prev: %h, now: %h -> STATE_PRECHARGE",
                                        activated_row_bank, active_addr[23:9]);
`endif
                        end
                    end else if (refresh_expired) begin
                        // Time to do a refresh.
                        sdram_cmd <= SDRAM_CMD_NOP;
                        sdram_dqm <= 2'b11;

                        auto_refresh_state_m <= STATE_AR_START;
                        state_m <= STATE_AUTO_REFRESH;
                    end else begin
                        sdram_cmd <= SDRAM_CMD_NOP;
                        sdram_dqm <= 2'b11;
                    end
                end

                STATE_READ_PENDING: begin
                    cas_latency <= {cas_latency[CAS_DELAY-1:0], 1'b0};
                    /*
                     * Read data appears on the DQ subject to the logic level on the DQM inputs two clocks earlier.
                     * If a given DQM signal was registered HIGH, the corresponding DQ will be High- Z two clocks later;
                     * if the DQM signal was registered LOW, the DQ will provide valid data (see ACTIVATE states).
                     */
                    sdram_cmd <= SDRAM_CMD_NOP;
                    if (cas_latency[CAS_DELAY]) begin
`ifdef D_SDRAM
                        $display($time, " SDRAM: STATE_READ_PENDING @[%h]: %h (next_word %h)", active_addr, sdram_d_i,
                                    next_word);
`endif
                        if (sel_i[3]) begin
                            if (next_word) begin
                                data_o[31:16] <= sdram_d_i;
                                sync_ack_o <= 1'b1;
                            end else begin
                                data_o[15:0] <= sdram_d_i;
                                transaction_start_q <= 1'b1;
                            end
                            next_word <= ~next_word;
                        end else begin
                            data_o <= sdram_d_i;
                            sync_ack_o <= 1'b1;
                        end
                        state_m <= STATE_ACTIVATED;
                    end else begin
                        sdram_dqm <= 2'b11;
                    end
                end

                STATE_PRECHARGE: begin
                    /*
                     * The PRECHARGE command is used to deactivate the open row in a particular bank or
                     * the open row in all banks. The bank(s) will be available for a subsequent
                     * row access a specified time (tRP) after the PRECHARGE command is issued.
                     */
                    precharge_all_task;

                    set_timer_task(TRP_CLKS);

                    state_m <= STATE_WAIT_TRP;
`ifdef D_SDRAM
                    $display($time, " SDRAM: STATE_PRECHARGE: -> STATE_WAIT_TRP");
`endif
                end

                STATE_WAIT_TRP: begin
                    if (timer_expired) begin
                        state_m <= STATE_IDLE;
`ifdef D_SDRAM
                        $display($time, " SDRAM: STATE_WAIT_TRP: -> STATE_IDLE");
`endif
                    end else begin
                        sdram_cmd <= SDRAM_CMD_NOP;
                    end
                end

                STATE_AUTO_REFRESH: begin
                    (* parallel_case, full_case *)
                    case (auto_refresh_state_m)
                        STATE_AR_START: begin
                            precharge_all_task;

                            set_timer_task(TRP_CLKS);

                            auto_refresh_state_m <= STATE_AR_WAIT_TRP;
                        end

                        STATE_AR_WAIT_TRP: begin
                            if (timer_expired) begin
                                sdram_cmd <= SDRAM_CMD_REFRESH;

                                set_timer_task(TRFC_CLKS);

                                auto_refresh_state_m <= STATE_AR_WAIT_TRFC;
                            end else begin
                                sdram_cmd <= SDRAM_CMD_NOP;
                            end
                        end

                        STATE_AR_WAIT_TRFC: begin
                            if (timer_expired) begin
                                reset_refresh_timer <= 1'b1;

                                state_m <= STATE_IDLE;
                            end else begin
                                sdram_cmd <= SDRAM_CMD_NOP;
                            end
                        end

                        default: begin
                            // Invalid state machine
                        end
                    endcase
                end

                default: begin
                    // Invalid state machine
                end
            endcase
        end
    end

endmodule
