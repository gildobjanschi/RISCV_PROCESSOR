/***********************************************************************************************************************
 * Copyright (c) 2024 Virgil Dobjanschi dobjanschivirgil@gmail.com
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy of this software and associated
 * documentation files (the "Software"), to deal in the Software without restriction, including without limitation the
 * rights to use, copy, modify, merge, publish, distribute, sublicense, and/or sell copies of the Software, and to
 * permit persons to whom the Software is furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in all copies or substantial portions of
 * the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE
 * WARRANTIES OF MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS
 * OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR
 * OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE SOFTWARE.
 **********************************************************************************************************************/

/***********************************************************************************************************************
 * This module implements an SPI master flash reader with a wishbone interface.
 *
 * It supports single and quad SPI (QPI) modes. If QPI_MODE is defined it will switch from SPI to QPI during reset
 * and it will operate in QPI mode after the module exists the reset state. Once it operates in QPI mode, to switch
 * back to SPI mode you need to restart the board. QPI -> SPI is not supported (nor very useful).
 *
 * The following datasheet applies: https://www.issi.com/WW/pdf/25LP-WP128F.pdf
 *
 * clk_i               -- The clock signal.
 * rst_i               -- Reset active high.
 * stb_i               -- The transaction starts on the posedge of this signal.
 * cyc_i               -- This signal is asserted for the duration of a cycle (same as stb_i).
 * addr_i              -- The address from where data is read
 * sel_i               -- The number of bytes to read (1 -> 4'b0001, 2 -> 4'b0011, 3 -> 4'b0111 or 4 bytes -> 4'b1111).
 * ack_o               -- The data request is complete on the posedge of this signal.
 * data_o              -- The data that was read (aligned to the least significant byte).
 * device_clk_i        -- Flash clock input generated by the PLL.
 * flash_csn           -- Flash chip select output.
 * flash_clk           -- Flash SPI clock output.
 * flash_mosi          -- Flash MOSI and QSPI bit 0.
 * flash_miso          -- Flash MISO and QSPI bit 1.
 * flash_wpn           -- Flash WP and QSPI bit 2.
 * flash_holdn         -- Flash HOLD and QSPI bit 3.
 **********************************************************************************************************************/
`timescale 1ns / 1ns
`default_nettype none

module flash_master #(parameter [31:0] FLASH_CLK_PERIOD_NS = 20) (
    // Wishbone interface
    input logic clk_i,
    input logic rst_i,
    input logic stb_i,
    input logic cyc_i,
    input logic [23:0] addr_i,
    input logic [3:0] sel_i,
    output logic ack_o,
    output logic [31:0] data_o,
    // The device clock is driving flash_clk
    input logic device_clk_i,
    // SPI flash wires
    output logic flash_csn,
    output logic flash_clk,
    inout logic flash_mosi,
    inout logic flash_miso,
    inout logic flash_wpn,
    inout logic flash_holdn);

    //==================================================================================================================
    // Flash device pin direction
    //==================================================================================================================
    logic qpi_mode = 1'b0;
    logic fpga_out_en = 1'b0;

    logic IO0_o = 1'b1, IO1_o = 1'b1, IO2_o = 1'b1, IO3_o = 1'b1;
    logic IO0_i, IO1_i, IO2_i, IO3_i;

    // In QPI mode flash_mosi, flash_wpn and flash_holdn are outputs (0) if fpga_out_en == 1.
    logic pin_0_2_3_dir;
    assign pin_0_2_3_dir = qpi_mode ? ~fpga_out_en : 1'b0;

    // In QPI mode flash_miso is an output (0) if fpga_out_en == 1.
    logic pin_1_dir;
    assign pin_1_dir = qpi_mode ? ~fpga_out_en : 1'b1;

    // .T = 0 -> pin is output; .T = 1 -> pin is input.
    TRELLIS_IO #(.DIR("BIDIR")) B0 (.B(flash_mosi), .I(IO0_o), .T(pin_0_2_3_dir), .O(IO0_i));
    TRELLIS_IO #(.DIR("BIDIR")) B1 (.B(flash_miso), .I(IO1_o), .T(pin_1_dir), .O(IO1_i));
    TRELLIS_IO #(.DIR("BIDIR")) B2 (.B(flash_wpn), .I(IO2_o), .T(pin_0_2_3_dir), .O(IO2_i));
    TRELLIS_IO #(.DIR("BIDIR")) B3 (.B(flash_holdn), .I(IO3_o), .T(pin_0_2_3_dir), .O(IO3_i));

    //==================================================================================================================
    // flash_clk drives the actual SPI flash clock and is enabled during SPI transactions.
    //==================================================================================================================
    logic clk_en = 1'b0;

    // Using the code below instead of: "assign flash_clk = clk_en ? device_clk_i : 1'b1;"
    // ensures that flash_clk will be initialized to 1'b1 at time = 0. Not doing so will trigger a flash_clk from
    // 0 -> 1 at time = 0 which starts a slave transaction (flash_csn = 0 at time = 0).
    logic man_flash_clk = 1'b1;
    assign flash_clk = clk_en ? device_clk_i : man_flash_clk;

    //==================================================================================================================
    // SPI state machine
    //==================================================================================================================
    // The state machine
    localparam [2:0] STATE_RESET = 3'b000;
    localparam [2:0] STATE_QPI_START = 3'b001;
    localparam [2:0] STATE_QPI_TX = 3'b010;
    localparam [2:0] STATE_QPI_DONE = 3'b011;
    localparam [2:0] STATE_IDLE = 3'b100;
    localparam [2:0] STATE_TX = 3'b101;
    localparam [2:0] STATE_RX = 3'b110;
    localparam [2:0] STATE_DONE = 3'b111;
    logic [2:0] state_m;

    // Rx and Tx buffers
    localparam SPI_BUFFER_SIZE = 32;
    logic [SPI_BUFFER_SIZE-1:0] spi_buffer;
    logic [31:0] spi_tx_clks, spi_rx_clks;
    logic [7:0] spi_dummy_clks;

    logic [2:0] reset_clks;

    logic sync_rst_i, sync_stb_i, sync_cyc_i;
    DFF_META dff_meta_rst (.reset(1'b0), .D(rst_i), .clk(clk_i), .Q(sync_rst_i));
    DFF_META dff_meta_stb (.reset(sync_rst_i), .D(stb_i), .clk(clk_i), .Q(sync_stb_i));
    DFF_META dff_meta_cyc (.reset(sync_rst_i), .D(cyc_i), .clk(clk_i), .Q(sync_cyc_i));

    //==================================================================================================================
    // Single wire TX SPI
    //==================================================================================================================
    task spi_tx_task(input [2:0] next_state_m);
        case (1'b1)
            |spi_tx_clks: begin
                clk_en <= 1'b1;
                /*
                * Data on the serial data lines need to be set tDS (Data In Setup Time) minimum 2ns before the
                * rising edge of flash_clk and needs to held for tDH (Data in Hold Time) minimum 2ns after the
				* rising edge of flash_clk.
                */
                IO0_o <= spi_buffer[31];
                spi_buffer[31:1] <= spi_buffer[30:0];

                spi_tx_clks <= {1'b0, spi_tx_clks[31:1]};
            end

            |spi_dummy_clks: begin
                spi_dummy_clks <= {1'b0, spi_dummy_clks[7:1]};
            end

            |spi_rx_clks: begin
                state_m <= STATE_RX;
            end

            default: begin
                clk_en <= 1'b0;
                /*
                    * flash_csn needs to be asserted tCH (CE# Hold Time) minimum 3ns after the rising edge of
                    * flash_clk used to send data on the serial line.
                    */
                flash_csn <= 1'b1;

                state_m <= next_state_m;
            end
        endcase
    endtask

`ifndef QPI_MODE
    //==================================================================================================================
    // Single wire RX SPI
    //==================================================================================================================
    task spi_rx_task(input [2:0] next_state_m);
        /*
         * The input data on the serial line is available after tV (Output Valid) maximum 5.5-7ns after the falling
         * edge of flash_clk. The time difference between the falling edge of flash_clk and the rising edge of clk_i
         * (used to read the data line) needs to be 7ns or greater.
         */
        spi_buffer <= {spi_buffer[SPI_BUFFER_SIZE-2 : 0], IO1_i};

        if (spi_rx_clks[0] == 1'b1) begin
`ifdef D_FLASH_MASTER_FINE
            $display($time, " FLASH_MASTER: Rx: %h", {spi_buffer[SPI_BUFFER_SIZE-2 : 0], IO1_i});
`endif
            clk_en <= 1'b0;
            /*
             * flash_csn needs to be asserted tCH (CE# Hold Time) minimum 3ns after the rising edge of
             * flash_clk used to send data on the serial line.
             */
            flash_csn <= 1'b1;

            state_m <= next_state_m;
        end else begin
            spi_rx_clks[30:0] <= spi_rx_clks[31:1];
        end
    endtask
`endif  // QPI_MODE

`ifdef QPI_MODE
    //==================================================================================================================
    // QUAD TX SPI
    //==================================================================================================================
    task qpi_tx_task(input [2:0] next_state_m);
        case (1'b1)
            |spi_tx_clks[7:0]: begin
                /*
                * Data on the serial data lines need to be set tDS (Data In Setup Time) minimum 2ns before the
                * rising edge of flash_clk and needs to held for tDH (Data in Hold Time) minimum 2ns after the rising
				* edge of flash_clk.
                */
                {IO3_o, IO2_o, IO1_o, IO0_o} <= spi_buffer[31:28];
                spi_buffer[31:4] <= spi_buffer[27:0];

                clk_en <= 1'b1;

                spi_tx_clks[7:0] <= {1'b0, spi_tx_clks[7:1]};
            end

            |spi_dummy_clks: begin
                fpga_out_en <= 1'b0;
                spi_dummy_clks <= {1'b0, spi_dummy_clks[7:1]};
            end

            |spi_rx_clks: begin
                fpga_out_en <= 1'b0;
                state_m <= STATE_RX;
            end

            default: begin
                fpga_out_en <= 1'b0;
                clk_en <= 1'b0;
                /*
                    * flash_csn needs to be asserted tCH (CE# Hold Time) minimum 3ns after the rising edge of
                    * flash_clk used to send data on the serial lines.
                    */
                flash_csn <= 1'b1;

                state_m <= next_state_m;
            end
        endcase
    endtask

    //==================================================================================================================
    // QUAD RX SPI
    //==================================================================================================================
    task qpi_rx_task(input [2:0] next_state_m);
        /*
         * The input data on the serial line is available after tV (Output Valid) maximum 5.5-7ns after the falling
         * edge of flash_clk. The time difference between the falling edge of flash_clk and the rising edge of clk_i
         * (used to read the data lines) needs to be 7ns or greater.
         */
        spi_buffer <= {spi_buffer[SPI_BUFFER_SIZE-5 : 0], IO3_i, IO2_i, IO1_i, IO0_i};

        if (spi_rx_clks[0] == 1'b1) begin
            clk_en <= 1'b0;
            /*
             * flash_csn needs to be asserted tCH (CE# Hold Time) minimum 3ns after the rising edge of
             * flash_clk used to send data on the serial lines.
             */
            flash_csn <= 1'b1;

            state_m <= next_state_m;
        end else begin
            spi_rx_clks[6:0] <= spi_rx_clks[7:1];
        end
    endtask

`endif  // QPI_MODE

    //==================================================================================================================
    // The SPI master
    //==================================================================================================================
    always @(posedge clk_i) begin
        if (sync_rst_i) begin
            clk_en <= 1'b0;

            fpga_out_en <= 1'b0;
            flash_csn <= 1'b1;
            ack_o <= 1'b0;

            reset_clks <= 3'b100;
            state_m <= STATE_RESET;
        end else begin
            if (ack_o) ack_o <= sync_stb_i;

            (* parallel_case, full_case *)
            case (state_m)
                STATE_RESET: begin
                    if (~|reset_clks) begin
                        flash_csn <= 1'b1;
`ifdef QPI_MODE
                        if (qpi_mode) begin
                            state_m <= STATE_IDLE;
                        end else begin
                            state_m <= STATE_QPI_START;
                        end
`else
                        state_m <= STATE_IDLE;
`endif
                    end else begin
                        flash_csn  <= 1'b0;
                        reset_clks <= {1'b0, reset_clks[2:1]};
                    end
                end

`ifdef QPI_MODE
                STATE_QPI_START: begin
`ifdef D_FLASH_MASTER
                    $display($time, " FLASH_MASTER: Entering QPI mode...");
`endif
                    // Send the command to switch to QPI
                    spi_buffer <= {8'h35, 24'b0};
                    spi_tx_clks <= 32'h0000_0080;

                    spi_rx_clks <= 32'h0000_0000;
                    spi_dummy_clks <= 8'h00;
                    /*
                    * tCS (CE# Setup Time) is the minimum time interval between the falling edge of flash_csn
                    * and the rising edge of the flash_clk. tCS = 3ns. flash_csn is asserted one clock cycle
                    * before the rising edge of flash_clk (which is enabled in the SPI tx/rx tasks).
                    */
                    flash_csn <= 1'b0;
                    state_m <= STATE_QPI_TX;
                end

                STATE_QPI_TX: begin
                    spi_tx_task(STATE_QPI_DONE);
                end

                STATE_QPI_DONE: begin
                    // Enter QPI mode
                    qpi_mode <= 1'b1;

                    state_m  <= STATE_IDLE;
`ifdef D_FLASH_MASTER
                    $display($time, " FLASH_MASTER: Entered QPI mode.");
`endif
                end
`endif  // QPI_MODE

                STATE_IDLE: begin
                    if (sync_stb_i & sync_cyc_i & ~ack_o) begin
`ifdef D_FLASH_MASTER_FINE
                        $display($time, " FLASH_MASTER: Read @[%h].", addr_i);
`endif
                        // Setup the Tx (command + 3 bytes of address) and the dummy cycles count
`ifdef QPI_MODE
                        spi_buffer <= {8'h0B, addr_i};
                        spi_dummy_clks <= 8'h20;  // 6 cycles
                        spi_tx_clks <= 32'h0000_0080;  // 8 nibbles

                        case (1'b1)
                            sel_i[3]: spi_rx_clks <= 32'h0000_0080;  // 8 nibbles
                            sel_i[1]: spi_rx_clks <= 32'h0000_0008;  // 4 nibbles
                            sel_i[0]: spi_rx_clks <= 32'h0000_0002;  // 2 nibbles
                            default:  spi_rx_clks <= 32'h0000_0002;  // 2 nibbles
                        endcase

                        fpga_out_en <= 1'b1;
`else  // QPI_MODE
                        if (FLASH_CLK_PERIOD_NS > 13) begin
                            // Normal read is more efficient (no dummy cycles) for flash_clk up to 80 MHz.
                            spi_buffer <= {8'h03, addr_i};
                            spi_dummy_clks <= 8'h00;  // 0 cycles
                        end else begin
                            // Fast read needs to be used for flash_clk > 80 MHz
                            spi_buffer <= {8'h0B, addr_i};
                            spi_dummy_clks <= 8'h80;  // 8 cycles
                        end
                        spi_tx_clks <= 32'h8000_0000;  // 32 bits

                        case (1'b1)
                            sel_i[3]: spi_rx_clks <= 32'h8000_0000;  // 32 bits
                            sel_i[1]: spi_rx_clks <= 32'h0000_8000;  // 16 bits
                            sel_i[0]: spi_rx_clks <= 32'h0000_0080;  // 8 bits
                            default:  spi_rx_clks <= 32'h0000_0080;  // 8 bits
                        endcase
`endif  // QPI_MODE
                        /*
                         * tCS (CE# Setup Time) is the minimum time interval between the falling edge of flash_csn
                         * and the rising edge of the flash_clk. tCS = 3ns. flash_csn is asserted one clock cycle
                         * before the rising edge of flash_clk (which is enabled in the SPI tx/rx tasks).
                         */
                        flash_csn <= 1'b0;

                        state_m   <= STATE_TX;
                    end
                end

                STATE_TX: begin
`ifdef QPI_MODE
                    qpi_tx_task(STATE_RX);
`else
                    spi_tx_task(STATE_RX);
`endif
                end

                STATE_RX: begin
`ifdef QPI_MODE
                    qpi_rx_task(STATE_DONE);
`else
                    spi_rx_task(STATE_DONE);
`endif
                end

                STATE_DONE: begin
                    // Data assembly for little endian
                    case (1'b1)
                        sel_i[3]: data_o <= {spi_buffer[7:0], spi_buffer[15:8], spi_buffer[23:16], spi_buffer[31:24]};
                        sel_i[1]: data_o[15:0] <= {spi_buffer[7:0], spi_buffer[15:8]};
                        sel_i[0]: data_o[7:0] <= spi_buffer[7:0];
                        default:  data_o <= 0;
                    endcase

                    ack_o   <= 1'b1;
                    state_m <= STATE_IDLE;
                end

                default: begin
                    state_m <= STATE_IDLE;  // This will never happen (invalid state machine)
                end
            endcase
        end
    end
endmodule
